.SUBCKT LED_red  K A
D1 1 A  LED_mod
V   K  1  DC 0
.MODEL LED_mod D (
+ IS=2.560e-014 N=3.007e+000 RS=8.513e-003
+ BV=6.100e+001 IBV=6.000e-006
+ EG=1.110e+000 XTI=3.000e+000
+ CJO=3.238e-011, M=3.388e-001 VJ=3.250e-001
+ FC=5.000e-001 KF=0.000e+000 AF=1.000e+000 )
.ENDS
