.subckt  seven_segmentda 1 2 3 4 5 6 7 8 10
V1 1a 1 DC 0
V2 2a 2 DC 0
V3 3a 3 DC 0
V4 4a 4 DC 0
V5 5a 5 DC 0
V6 6a 6 DC 0
V7 7a 7 DC 0
V8 8a 8 DC 0
D1 10 1a DLEDSEG
D2 10 2a DLEDSEG
D3 10 3a DLEDSEG
D4 10 4a DLEDSEG
D5 10 5a DLEDSEG
D6 10 6a DLEDSEG
D7 10 7a DLEDSEG
D8 10 8a DLEDSEG
.MODEL DLEDSEG  D (
+ IS=2.560e-014 N=3.007e+000 RS=8.513e-003
+ BV=6.100e+001 IBV=6.000e-006
+ EG=1.110e+000 XTI=3.000e+000 
+ CJO=3.238e-011, M=3.388e-001 VJ=3.250e-001
+ FC=5.000e-001 KF=0.000e+000 AF=1.000e+000 )
.ends