*2N6426 MCE 6/19/97
*Ref: Motorola Small-Signal Device Databook, Q4/94
*Si 625mW 40V 500mA pkg:TO-92B 1,2,3
.SUBCKT 2N6426   1 2 3
*    TERMINALS:  C B E
Q1 1 2 4 QPWR .1
Q2 1 4 3 QPWR
.MODEL QPWR NPN (IS=600F NF=1 BF=368 VAF=114 IKF=0.4 ISE=13.3P NE=2
+ BR=4 NR=1 VAR=48 IKR=0.6 RE=0.2 RB=0.8 RC=80M CJE=147P XTB=1.5
+ VJE=0.74 MJE=0.45 CJC=9.4P VJC=1.1 MJC=0.24 TF=69.6N TR=3.01U)
.ENDS 
* Origin: Mcebjt.lib
