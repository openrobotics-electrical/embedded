**************** Power Discrete MOSFET Electrical Circuit Model *****************
* Product Name: FQP7P06
* 60V P-Channel MOSFET and TO-220* Creation : Nov.-04-2002 * Fairchild Semiconductor
*--------------------------------------------------------------------------------
.SUBCKT FQP7P06 20 10 30
Rg 10 1  1
M1 2 1 3 3 DMOS  L=1U  W=1U
.MODEL DMOS PMOS (VTO={-3.00*{-0.00048*TEMP+1.012}} KP={4*{-0.00046*TEMP+1.0115}}
+ THETA=0.056  VMAX=1.30E5   LEVEL=3)
Cgs 1 3 200P
Rd 20 4 0.1  TC=0.007
Dds 4 3 DDS
.MODEL DDS D(BV={60*{0.0011*TEMP+0.9725}}  M=0.37   CJO=85P   VJ=0.609)
Dbody 20 3 DBODY
.MODEL DBODY D(IS=3.0E-13  N=1.0  RS=0.0012  EG=1.15  TT=77n)
Ra 4 2  0.1  TC=0.007
Rs 3 5  0.075
Ls 5 30 5n
M2 1 8 6 6 INTER
E2 8 6 4 1 2
.MODEL INTER PMOS (VTO=0 KP=10 LEVEL=1)
Cgdmax 7 4 330P
Rcgd 7 4 1E7
Dgd  4 6 DGD
Rdgd 4 6 1E7
.MODEL DGD D(M=0.54 CJO=330P VJ=0.52)
M3 7 9 1 1 INTER
E3 9 1 4 1 -2
.ENDS FQP7P06